function Bit#(32) shiftRightPow2(Bit#(1) en, Bit#(32) unshifted, Integer power);
    return 0;
endfunction

function Bit#(32) barrelShifterRight(Bit#(32) in, Bit#(5) shiftBy);
    return 0;
endfunction